-- IndividualPWMLEDController.vhd
-- 2025.03.23
--
-- Takes in PWM cycle data and controls an LED's brightness
-- TODO: find a better file and entity name
-- TODO: add state selector so "set brghtness", "increase brightness", etc.
-- Maybe implement gamma correction in this component

library ieee;
library lpm;

use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use lpm.lpm_components.all;

entity singleledcontroller is
port(
    latch       : in  std_logic; -- Latches cycle data to saved state when 1
    input_cycles : in  integer;   -- Number of clock ticks you want the led to be on
    total_cycles: in  integer;   -- Total number of clock ticks total for one PWM period
    clock       : in  std_logic; -- Referenced for PWM brightness
    led_out     : out std_logic  -- Physical output for a singular LED
    );
end singleledcontroller;

architecture a of singleledcontroller is
    signal total_count  : integer; -- Total amount of clock cycles in one PWM period minus 1 so input 1023 for 1024 total cycles
    signal on_count     : integer; -- Amount of clock cycles where LED is on
    signal ticks        : integer := 0; -- Counter to determine LED state if counter <= on_count LED is on else LED is off
begin
    
    process (latch, clock)
    begin
        if (latch = '1') then -- latch necessary values
            total_count <= total_cycles; 
            on_count <= input_cycles;
        end if;
        if (rising_edge(clock)) then
			ticks <= ticks + 1;
        end if;
        if (ticks > total_count) then
            ticks <= 0;
        end if;
    end process;

    led_out <= '1' when (ticks < on_count) else '0';
end a;
